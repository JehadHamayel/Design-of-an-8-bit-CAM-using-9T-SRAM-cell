*** SPICE deck for cell nand{sch} from library Project
*** Created on Sat Jun 24, 2023 14:15:13
*** Last revised on Thu Jul 06, 2023 08:45:54
*** Written on Thu Jul 06, 2023 08:49:50 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: nand{sch}
Mnmos@8 out h net@79 gnd NMOS L=0.044U W=0.22U
Mnmos@9 net@79 g net@80 gnd NMOS L=0.044U W=0.22U
Mnmos@10 net@80 f net@81 gnd NMOS L=0.044U W=0.22U
Mnmos@11 net@81 e net@82 gnd NMOS L=0.044U W=0.22U
Mnmos@12 net@82 d net@83 gnd NMOS L=0.044U W=0.22U
Mnmos@13 net@83 c net@84 gnd NMOS L=0.044U W=0.22U
Mnmos@14 net@84 b net@86 gnd NMOS L=0.044U W=0.22U
Mnmos@15 net@86 a gnd gnd NMOS L=0.044U W=0.22U
Mpmos@0 vdd h out vdd PMOS L=0.044U W=0.22U
Mpmos@1 vdd g out vdd PMOS L=0.044U W=0.22U
Mpmos@2 vdd f out vdd PMOS L=0.044U W=0.22U
Mpmos@3 vdd e out vdd PMOS L=0.044U W=0.22U
Mpmos@4 vdd d out vdd PMOS L=0.044U W=0.22U
Mpmos@5 vdd c out vdd PMOS L=0.044U W=0.22U
Mpmos@6 vdd b out vdd PMOS L=0.044U W=0.22U
Mpmos@7 vdd a out vdd PMOS L=0.044U W=0.22U

* Spice Code nodes in cell cell 'nand{sch}'
vdd vdd 0 dc 1.3
va a 0 pulse 1.3 0 1p 1p 1p 150n 300n
vb b 0 pulse 1.3 0 1p 1p 1p 300n 600n
vc c 0 pulse 1.3 0 1p 1p 1p 600n 1200n
vd d 0 pulse 1.3 0 1p 1p 1p 1200n 2400n
ve e 0 pulse 1.3 0 1p 1p 1p 2400n 4800n
vf f 0 pulse 1.3 0 1p 1p 1p 4800n 9600n
vg g 0 pulse 1.3 0 1p 1p 1p 9600n 19200n
vh h 0 pulse 1.3 0 1p 1p 1p 19200n 38400n
cload out 0 200fF
.tran 76800n 
.include C:\elec\22nm.txt
.END
